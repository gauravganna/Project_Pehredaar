--VHDL code for 4 Digit BCD Counter created by Gaurav Ganna as part of Project Pehredar
--Date 29/03/2018
library ieee;							-- Library Declaration
use ieee.std_logic_1164.all;		-- Use std_logic_1164 package from ieee library
use work.RFID_Project.all;			-- Include the package created as part of Project

entity DGT_4_Counter is
	port(
	);